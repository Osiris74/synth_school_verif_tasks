`timescale 1ns/100ps

module testbench;

    logic [31:0] A;
    logic [31:0] B;
    logic [31:0] C;

    logic [7:0] increment;

    sum DUT(
        .a ( A ),
        .b ( B ),
        .c ( C )
    );

    `include "checker.svh"

    initial begin

        // TODO:
        // Представьте, что для каждого входного операнда (A и B)
        // интервал всех возможных значений равномерно разбит на
        // 8 одинаковых по размеру подинтервалов:
        
        // |0....|.....|.....|.....|.....|.....|.....|..max|
        // |  0  |  1  |  2  |  3  |  4  |  5  |  6  |  7  |
    
        // Ваша задача - подать значения из каждого интервала для
        // каждого операнда.
        
        // В конце симуляции будет выведена статистика о том, какая
        // часть из требуемых значений была подана. Для оценки того,
        // значения из какого интервала не были поданы, воспользуйтесь
        // отчетом 01_sum/stats/covsummary.html (отчет сформируется
        // после завершения симуляции).

        // Не забудьте про выставление задержек через '#'!

        // Пишите внутри этого блока
        //------------------------------------------------------------
        increment = 255;

        for (int i=0; i<increment; i++) 
        begin
          #10; A [7:0]   = i; B[7:0]   = i; 
          #10; A [15:8]  = i; B[15:8]  = i;
          #10; A [23:16] = i; B[23:16] = i;   
          #10; A [31:24] = i; B[31:24] = i;
        end 
        //------------------------------------------------------------

        -> gen_done;

    end

endmodule
